module fv_tb;

  arbiter_sva #(4) inst1();

  arbiter_sva #(7) inst2();

endmodule
